library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity secded_test_32bits is
	port( address : in std_logic_vector(10 downto 0);
		clk : in std_logic;
		dout : out std_logic_vector(42 downto 0));
	end;

architecture v1 of secded_test_32bits is

	constant ROM_WIDTH: INTEGER:= 43;
	constant ROM_LENGTH: INTEGER:= 2048;

	subtype rom_word is std_logic_vector(ROM_WIDTH-1 downto 0);
	type rom_table is array (0 to ROM_LENGTH-1) of rom_word;

constant rom: rom_table := rom_table'(
	"0111100000000000000000000000000000000000000",
	"0110110000000000000000000000000000001000101",
	"0110110000000000000000000000000000000000100",
	"0110100000000000000000000000000000000000001",
	"0100000001000000000000000000000000001011110",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010000",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010010",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010011",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010100",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010101",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010110",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010111",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011000",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011001",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011010",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011011",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011100",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011101",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001010001",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000001000101",
	"0100000001000000000000000000000000001011111",
	"0010000011000010000000000000000000000000000",
	"0110110000000000000000000000000000001101101",
	"0110110000000000000000000000000000010000001",
	"0100100000000000000000000000000000000000000",
	"0100000001000000000000000000001000100010001",
	"0000010001000000000000000000000000010000000",
	"0110100010100000000000000000000000001000101",
	"0110110000000000000000000000000000001100110",
	"0000000001100000000000000000000000000001001",
	"0110110000000000000000000000000000001011111",
	"0101000001000000000000000000000000000001110",
	"0100000000000000000000000000001000100010001",
	"0000010000000000000000000000000000010000000",
	"0010100001000000000000000000000000000000000",
	"0001100001100000000000000000000000000000001",
	"0110100010100000000000000000000000001001010",
	"0100100000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0100010000000000000000000000001000100010001",
	"0110110000000000000000000000000000001011111",
	"0000000001100000000000000000000000000001000",
	"0100010000100000000000000000001000100010001",
	"0110110000000000000000000000000000001011111",
	"0101000000100000000000000000000000000001110",
	"0001100001100000000000000000000000000000001",
	"0110100010100000000000000000000000001010110",
	"0000000000000000000000000000000000011111111",
	"0100010000000000000000000000001000100010001",
	"0110110000000000000000000000000000001011111",
	"0100100000000000000000000000000000000000000",
	"0000000010000000000000000000000000000000001",
	"0000000010100000000000000000000000011010110",
	"0001100010100000000000000000000000000000001",
	"0110100010100000000000000000000000001100001",
	"0001100010000000000000000000000000000000001",
	"0110100010100000000000000000000000001100000",
	"0100100000000000000000000000000000000000000",
	"0000000010000000000000000000000000000000010",
	"0000000010100000000000000000000000000110100",
	"0001100010100000000000000000000000000000001",
	"0110100010100000000000000000000000001101000",
	"0001100010000000000000000000000000000000001",
	"0110100010100000000000000000000000001100111",
	"0100100000000000000000000000000000000000000",
	"0000000011100000000000000000000000000100000",
	"0010000100000110000000000000000000000000000",
	"0000010100010000000000000000000000000000000",
	"0000100100000000000000000000000000000000000",
	"0110100010100000000000000000000000001111011",
	"0110100000000000000000000000000000001111110",
	"0101000011000000000000000000000000000000100",
	"0001100011100000000000000000000000000000001",
	"0110100010100000000000000000000000001101110",
	"0000000000100000000000000000000000000001010",
	"0110110000000000000000000000000000001010010",
	"0000000000100000000000000000000000000001101",
	"0110110000000000000000000000000000001010010",
	"0100100000000000000000000000000000000000000",
	"0000000000100000000000000000000000000110001",
	"0110110000000000000000000000000000001010010",
	"0110100000000000000000000000000000001110011",
	"0000000000100000000000000000000000000110000",
	"0110110000000000000000000000000000001010010",
	"0110100000000000000000000000000000001110011",
	"0000000000100000000000000000000000000001010",
	"0110110000000000000000000000000000001010010",
	"0000000000100000000000000000000000000001101",
	"0110110000000000000000000000000000001010010",
	"0100100000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000");

begin

process (clk)
begin
	if clk'event and clk = '1' then
		dout <= rom(conv_integer(address));
	end if;
end process;
end v1;
